// Example 4 - incomplete rn
module four-bit-shift-register (
    input wire i_clk,
    input reg [3:0]
);
    begin
    end
endmodule